module PCTarget (
    input  logic [31:0] PCE,
    input  logic [31:0] ImmExtE,
    output logic [31:0] PCTargetE
);
    always_comb begin
        PCTargetE = PCE + ImmExtE;
    end
endmodule
